module control_tb();
  
  reg clock;
  
  control_unit_data_processing datapath1(clock);
  
  initial
  begin
  clock=0;
  end
  
  always
  begin
  #10 clock=~clock;
  end
  
endmodule
