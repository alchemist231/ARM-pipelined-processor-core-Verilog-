module instantiate_tb();
  register_file_tb trial();
  
endmodule
