module and_tb();
  wire c;
  reg a,b;
  
  and1 a1(a,b,c);
  
  initial 
  begin
    a=0;  b=0;
 
 end
 endmodule
 