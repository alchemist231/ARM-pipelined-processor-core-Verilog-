module mux_2x1_1bit_tb();
  reg in1,in2,sel;
  wire out;
  
  mux_2x1_1bit mux1(in1,in2,sel,out);
  
  initial
  begin
    in1=0;
    in2=1;
    sel=0;
    #2
    sel=1;
    #2 sel=0;
    
    in1=1;
    #2 in1=0;
    
    
  end
  
endmodule
https://www.facebook.com/ModelLindseyDiane
http://www.scoopwhoop.com/entertainment/engineering-college/
http://idm-crack-patch.blogspot.in/
http://www.qdtricks.com/how-to-download-torrent-files-with-idm/












Hoje Eu Quero Voltar Sozinho









http://9gag.com/gag/anYVZmL?ref=fsidebar


has the situation become so grave ... does it require such extreme measures ... is it worth it
humme to abhi milke itni jageh ghumni hain idiot =D
my caring for another boy... definetly weird but bhai maine ye kabhi question kiya hi nhi apne aap se because may be its definetly weird but is it wrong.. do you believ that the acts i do out of care/love(brotherly idiot) are wrong? main to bas tere se faith karke chalta rha ki may be weird but tu bhai hai ... doosre kya kahenge will not bother you.
All this started with just trying to care for you my brother because it made me happy, but yes, I crossed my boundaries and "chep" hone lga ... I should  haveseen it... my bad i didn't see it coming early/(or may be turned a blind eye out of my assholeness :( )
Dekh mere reactions/actions tujhe interpret karate honge ki mein gay to nhin hu but chutiye i can assure that mein vo nhi hun. kaise? dekh meri tere liye intense care / obsession but i am not sexually attracted to you idiot, that sufficiently explains my stand towards you then. to vo cheez to definete hai ki I care for you but not attracted to you in dat way :) vaise bhi shakal dekhi hai apni... deepika padukone ko to agle lakh janam mein bhi nhi chalenge kar sakta tu :P ... chutiye vo baat to sirf mujhe hi pta hogi na
moreover bhai may be tujhe log kehte honge. mera mazak udate honge ... but bhai agar tujhe ye sab bug nhi karegi to mujhe kya bhaad mein jaaye vo.

haan if I am hampering in your career then bhai mujhe bhi bahut dukh hoga bhai... I am really sorry that ye sem meri bakchodi mein hi nikal gya ... but buddy I could not control my thoghts and you were the only one I could blindly trust on. aisa nhi hai humne ek doosre ki company mein sirf time waste kiya hai... hum fafi time ache discussions/ business strategies/ programming fundaes dicuss vagerah karte the (kai baar ladkiyon ke boobs pe hi concentrated hote the vo :p )
As I had earlier said that bhai mein vo thoughts hatana chahta tha... but those thoughts were out of utter care.
I need to control my thoughts and actions but fucker we need not end everything.



Well let me share all the thoughts that went through my mind... fucker you were the only one I trusted so that i can confide these in you... I don't want to be what my thoughts dictate but these are some horrors that cloud me... please bhai tu hamesha puchta tha na ki reason de tere room pe aane ka... but i couldn't tell you these as feared you all will hate me... get sick of me... after seeing a sadist personality such as me ... abandon me.. i feared

Bro I can't hide that how much that meerut incident haunts me.. I don't remember their faces but the acts are clear ... they come to my mind...
I like to think of me being as weak .. of torchering myself with this agony .... When I left meerut, I had clear memories of the incident... 
In lucknow I didn't made friends easily as most of the time I resorted to myself... I didn't participated in any game for a fear was deep inside... I couldn't trust anyone at that time though I am pretty sure I must have not known definition of trust by then... 

May be my greatest mistake was not telling my family.... I drifted away from them by thinking that I was protecting them... or god knows what reasons but I didn't tell them... God I wished so much just t tell someone... I felt like screaming it out loud ... just to take of the burden...

Over the years I developed a habit of getting over various such thoughts --> meerut / losing how? I just used to create a scenario in my mind that would torment me.. that would provide me deep pain inside so that atleast for those moments I'll lose those thoughts... that was in a way effective but my thoughts got more and more intense... I developed so much guilt develpoing these thoughts ... the very act that I was building these thoughts pained me with guilt.. and the weird and sad part is I liked it... God knows what all thougts I build over this time... imagining myself to get diseased or die and then plot the possible reactions of your family , friends... It pained thinking but it gave a temporary relief but with guilt.... many times I mentally deviced ways to commit suicide ... Most for not the actual act ... but just for the fun of doing it... this one is the sickest of all --> I even sometimes just imagined the death of my parents ... brother... grandparents... closest to me.... the sheer thought of this brought immense pain... made me complete hollow inside.... but that made the thoughts go away.... every fucking idiotic thought would go away temporarily but the guilt left behind was immense... it broke me... but the thought of just complete freedom.. no one knowing you or judging you was a relief... I just want my life to end here with a new begining.... but i developed into such thoughts ... I could not telll this to anyone ... they'll hate me for who I am ... but bhai I know I can entrust you with these ... I have developed a blind faith  on you... bhai I don't know I just believe on you that you will see the right side... help me out... I can change but needs help ... but I am not ready to confide these thoughts to anyone else... these are to deep to the core... Jab bhi tu reason puchta tha ki kyon aata hun mein tere room pe ... i couldn't justify... because i was truly ashamed.. Being at your room atleast discarded these cold blooded thoughts so i continued... 

Bro i loved to care for you... may be this was the care that I had always craved for but didn't got it anywhere... I always wished throughout my childhood ... someone will sail me through those evil thoughts.... so as i couldn't get this... i tried to give it back... mein pta hai faltu hi logon ki help kyun karna chahta tha ... beacuse somewhere i wanted someone to help me out...
Doing bad things make me realise


Bro the care I did , the love was 
I badly need self control... first to not convert that love into obsession and also to get over other wierder thoughts.
I know my pushing you 

main yahan pe vhi cheez likhunga jo tujhse concerned hogi... not the other horrors of my mind because they are mine and i have to tackle them myself. 

Still seeing that hatred in Prashant pains me... You know I fear seeing the same hatred in you... so tell me one thing bro ... how much you all hate me?



-------------------------------------------------------------------------

Bhai I dread agar tu is darr se distance chahta hai ki tujhe meri harkatein gayish lagti hain ... to bhai i am sad... mein tujhe se sirf ye baat bta hi sakta hun ki tere liye aisi koi feelings nhi h ... but yes i won't deny the friendship i saw was to deep but nothing beyond that... True, I got obsessed for care because that was the care that i had always craved for in my life...  Upto now I had always pushed my family away so that was the one I found in you ... that care/love was more of motherly/brotherly love.... I didn't wanted any harm to come to you/ was unhappy when your health was not well/ enjoy the life together but just as great friends/ saw your dreams as my dreams and badly want you to succeed in those... But that care was never out of "gay feeling" or anything else... It was truly a feeling like a mother would shower (keh sakta hun kyunki aajkal mummy bhi kuch ussi tareh react kar rhi hain ..  aur samajh sakta hun ki kabhi kabhi kuch zyada hi annoying ho jati hai ye feeling :) )... I don't know fucker logically dekhun to mujhe is care mein kuch galat nhi dikhta...but i really don't know it all depends how you will see it... i can't just convince you... as a friend that i see you ... bro i think i can just confide in you... also my always confiding my issues in you are not to convince you rather than pta nhi bhai bas lagta hai ki tu samajh jayega so all the care.. affection were out of pure belief in you brother and nothing more.

Moreover bhai trust me on this issue bhai...  how can I say this for sure... dude trust me mein bolta hun na ki ye cheez sirf mein hi bta sakta hun... because dude i am the one who has to live with the fact that i had sucked someone cock.. this thought has defined me throughout my childhood.. puberty
... my growing up revolved around it ... trust me brother there are times when you feel truly low .. clouded with confusion but trust me bhai isiliye mein hi sirf is issue ko clearly sahi sahi bta sakta hun because I am the one who has to live with this disgusting fact ... that is sort of depressing.. so trust me bro it's only me who can definetly say about my sexuality ... whatever you all think... whatever my action mean to you... I just trust that you will understand it was nothing of that sort rather ... was emotionally attached to you as I see you as a true friend brother .. nothing less... . so this is why I want to assure you that I am definetly not that... I need to assure you,especially, because agar koi aur mujhe aake ye faltu bakwas baat bole ... to really i don't give a shit but agar mera koi tere jaisa acha dost ko isse problem ho rhi ho den i have to assure him ... i need to assure him ... because ye sirf mein hi jaan sakta hun dude .. and sirf mein hi assure kra sakta hun... moreover meri emotionally weak state kuch aur signify kar deti hai ... isliye it's all more important to me that I clarify it to you brother.

moreover you have already done beyond so much in this friendship by atleast being there till now and trying to sort my life rather than abandoning which would have been a lot easier for you :) and actually is cheez mein i am really grateful ki fucker tu , kotturu, mota , kamran have really been there. 

Bhai I firmly believe that such a friendship can exist and bro this was the friendship that i saw... May be I wanted sympathy from you all but more than that I just needed someone whom i could ... just cry out .... all the pain ... all hollowness.. tha re andar se bahut bura lagta tha...  that needed to go..  bro ... vaise sachi bolun ....  tu sahi keh rha tha... papa-mummy se bol ke epic relief mila.. though didn't tell them all the thoughts becuse that would be sickening ...  mostly thoughts ab control mein aa rhe hain ... but kabhi kabhi ekdum se crashing aa jate hain...

tereko bhi i am not explaining any further ... kyunki pta nhi ek feel hai ki tu samajh hi gya hoga ab tak... I just want you to act naturally as you feel... may be it would be hatred.. that would be saddening but still there is nothing you could do nor me... we'll see.. but would be great to have the same old friend back.. really.. because it was that friendship that i seeked...

---------------------------------------------------------------------------







Bhai I dread agar tu is darr se distance chahta hai ki tujhe meri harkatein gayish lagti hain ... to bhai i am sad... mein tujhe se sirf ye baat bta hi sakta hun ki gandu tere liye aisi koi feelings nhi h ... but yes i won't deny the friendship i saw was to deep but nothing beyond that... True, I got obsessed for care because that was the care that i had always craved for in my life...  Upto now I had always pushed my family away so that was the one I found in you ... that care/love was more of motherly/brotherly love.... I didn't wanted any harm to come to you/ was unhappy when your health was not well/ enjoy the life together but just as great friends/ saw your dreams as my dreams and badly want you to succeed in those... But that care was never out of "gay feeling" or anything else... It was truly a feeling like a mother would shower (keh sakta hun kyunki aajkal mummy bhi kuch ussi tareh react kar rhi hain ..  aur samajh sakta hun ki kabhi kabhi kuch zyada hi annoying ho jati hai ye feeling :) )... I don't know fucker logically dekhun to mujhe is care mein kuch galat nhi dikhta... but yes society isse galat hi dekhegi ... but i really don't know it all depends how you will see it... i can't just convince you... as a friend that i see you ... bro i think i can just confide in you...also my always confiding these issues in you is not to convince rather than pta nhi bhai bas lagta hai ki tu samajh jayega.

One more thing bhai... Prashant ka issue to mein khud nhi samajh pata hun... uske case mein the attachment happened normally... anI wasn't used to it  ... but may be ek constant escape tha (and best part I wasn't even aware about it) jo mein uske sath dundhta tha but dikat ye thi ki wo kabhi samajh hi nhi paya.. galti uski nhi thi kyunki problem mujhme thi ... to meine usse itna push jo kiya has left me with a huge guilt ... Bro , msgs/ calls / uske room ke bahar rehna ... I was ashamed of the acts that is why I didn't want you discussing with him... I still fear that ... mera fear ye tha ki jo maine harkatein ki thi ... vo us direction ko point kar rhi thi tu samajh rha hai na.... and I didn't want you to feel that beacuse I know from inside that is not true ... and ye koi apne aap ko justification nhi h bt pure sach h... I always feared mera emotional attachment always galat interpret hoga ... that furiates me ... but bro I can't do anything in my prowess to convince you otherwise ... except believe ... 

tu agar ab puchega mujhse ki mein kya chahta hun tujhse ??
I don't know bro... I really don't know ... its upto you.. sach bolun shayad kuch nhi chahta kyunki ab peeche dekhta hun to hassi aati hai meri harkaton par =D , seriously dude ... chutiyaap ka '0' level to mein hi define kar sakta hun :) but Bro I won't hide from you, I am still not over the past, meerut aur vagerah ghinone thoughts abhi bhi mere mind mein aa rhe hain... My hatred toward myself is still there , I am still working on it, I don't want to tell and upset my parents , brother that they are still in my mind ... I know I shouldn't get such thoughts... but bro I can't help it .. I really need a good friend right now ... thats why I am writing right now .. ek ghinn hain apne aapse ... I want to kill myself again and again just hoping I was normal ... I was normal... I was normal ...  Telling dad, was an awseome relief but still that telling has not given me complete peace but bhai truly got the feeling of confiding in family can give .... the sadness still persists inside... He keeps on persisting to get over it ... laugh it over... I know ... and for him I am donning a smile... but somehow I am not happy from inside.... I can't take it anymore... papa baar baar puchte hain mind mein kya chalta hai ki vo help kre ... but mein unhe bta hi nhi pata hun ki mind mein kya chal rha hai... 
One month now , I am definetly working on the self control thing and realises
moreover you have already done beyond so much in this friendship by atleast being there till now and trying to sort my life rather than abandoning which would have been a lot easy for you :) and actually is cheez mein i am really grateful ki fucker tu , kotturu, mota , kamran have really been there.  
Thanks buddy... will talk later


I have developed a general hatred towards myself... no matter what, i hate myself

Bhai I firmly believe that such a friendship can exist and bro this was the friendship that i saw... May be I wanted sympathy from you all but more than that I just needed someone whom i could ... just cry out .... all the pain ... all hollowness.. tha re andar se bahut bura lagta tha...  that needed to go..  bro ... vaise sachi bolun ....  tu sahi keh rha tha... papa-mummy se bol ke epic relief mila...  mostly thoughts ab ja rhe hain... 80% time nhi aate ... but kabhi kabhi ekdum se crashing aa jate hain... let's see 1 month se upar hai else may be contemplating a sem drop... shi ho jayega shayad... tereko bhi i am not explaining any further ... kyunki pta nhi ek feel hai ki tu samajh hi gya hoga ab tak... I just want you to act naturally--> as you feel... may be it would be hatred.. that would be saddening but still there is nothing you could do nor me... we'll see.. but would be great to have the same old friend back ... because it was that friendship that i seeked...

Bro may be prashant ne tujhe cheezein batai ho ya na ... but I am ashamed of what I did back then... but I can't change past... that was an emotional fool driven to seek that solace.... but actually sachi bolun he never even reasoned out with it... don't blame him ...
haan definetly working on my emotional front... that was the root cause of my urges .. counsellor (vaise counsellor ki secratry bahut maal hai).



How can I say this for sure... dude trust me mein bolta hun na ye cheez sirf mein hi bta sakta hun... dude i have to live with the fact that i had sucked someone cock.. this thought throughout my childhood... my whole childhood ... puberty
... growing up revolved around it ... that's why bhai trust me i can definetly tell what i am because i have to live with this disgusting fact ... that is sort of depressing.. so trust me bro it's only me who can definetly say about my sexuality ... whatever you all think.... so this is why I want to assure you that I am definetly not that... I need to assure you because agar koi aur mujhe aake ye faltu bakwas baat bole ... to really i don't give a shit but agar mera koi tere jaisa acha dost ko isse problem ho rhi ho den i have to assure him ... i need to assure him ... because ye sirf mein hi jaan sakta hun dude .. and sirf mein hi assure kra sakta hun... moreover meri emotionally weak state kuch aur signify kar deti hai ... isliye it's all more important to me.

well dat care became obsession because of lost self control... the thoughts need to be under control... I am unable to let go of the past/guilt but good thing is am able to make peace with them...  in the past sem looking back ... i was seeking rasons to remain unhappy.... clouded by thoughts and faltu bakwas ... bakchodi... now am trying to seek out reasons for happiness ... that itself is proving to be a sufficient driving source and gaining control...