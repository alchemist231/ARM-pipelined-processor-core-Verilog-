module pc_incrementer(pc_current,pc_increment,pc_next);
  input [31:0] pc_current;
  input pc_increment;
  output [31:0] pc_next;
  
  wire [31:0] pc_current;
  wire pc_increment;
  wire [31:0] pc_next;
  
  //later include exception handling if overflow in pc address????
  
  assign pc_next=(pc_increment==1)? pc_current+4:pc_next;
  
endmodule
