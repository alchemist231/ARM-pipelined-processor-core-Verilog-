module shifter(enable,in_data,in_data_imm,imm_or_reg,shift_control,shift_amt_imm,shift_amt_reg,rotation_code,carry_in,carry_out,out_data);
  
  input [31:0] in_data,shift_amt_reg;
  input enable,carry_in,imm_or_reg;
  input [7:0] in_data_imm;
  input [3:0] rotation_code;
  input [4:0] shift_amt_imm;
  input [2:0] shift_control;
  
  output [31:0] out_data;
  output carry_out;
  
  wire [31:0] in_data,shift_amt_reg;
  wire [7:0] in_data_imm;
  wire [2:0] shift_control;
  wire [4:0] shift_amt_imm;
  wire enable,carry_in,imm_or_reg;
  reg sign_bit;
  reg [31:0] out_data;
  reg carry_out;
  
  reg [4:0] temp;
  reg [31:0] temp1;
  
  initial
  begin
  out_data=32'h0;
  carry_out=0;
  end
  
  
  always@(enable,in_data,in_data_imm,imm_or_reg,shift_control,shift_amt_imm,shift_amt_reg,rotation_code,carry_in)
  begin
    if(enable)
      begin
      if(~imm_or_reg)
      begin
      case(shift_control)
        3'b000 :begin
                if(shift_amt_imm!=0)
                  begin
                    carry_out=in_data[31-shift_amt_imm+1];
                    out_data=in_data<<shift_amt_imm;
                  end
                else
                  begin
                    carry_out=carry_in;
                    out_data=in_data;
                  end
                end
                
        3'b001 :begin
                if(shift_amt_reg!=0)
                  begin
                    carry_out=in_data[31-shift_amt_reg+1];
                    out_data=in_data<<shift_amt_reg;
                  end
                else
                 begin
                    carry_out=carry_in;
                    out_data=in_data;
                 end
                end
                
        3'b010 :begin
                if(shift_amt_imm!=0)
                  begin
                    carry_out=in_data[shift_amt_imm-1];
                    out_data=in_data>>shift_amt_imm;
                  end
                else
                 begin
                   carry_out=carry_in;
                  out_data=in_data;
                 end
                end
                
        3'b011 :begin
                out_data=in_data>>shift_amt_reg;
                if(shift_amt_reg!=0)
                    carry_out=in_data[shift_amt_reg-1];
                else
                    carry_out=carry_out;
                end
                
        3'b100 :begin
                sign_bit=in_data[31];
                temp=shift_amt_imm;
                out_data=in_data;
                while(temp>0)
                begin
                  out_data={sign_bit,out_data[31:1]};
                  temp=temp-1;
                end
                // out_data={sign_bit[shift_amt_imm-1:0],in_data[31:shift_amt_imm]};
                if(shift_amt_imm)
                    carry_out=in_data[shift_amt_imm-1];
                else
                    carry_out=carry_out;
                end
                
       3'b101 :begin
               if(|shift_amt_reg[31:5])
                  begin
                  out_data={32{in_data[31]}}; 
                  carry_out=1; 
                  end              
               else
                 sign_bit=in_data[31];
                 out_data=in_data;
                 temp1=shift_amt_reg;
                 while(temp1!=0)
                 begin
                   out_data={sign_bit,out_data[31:1]};
                   temp=temp-1;
                 end
              //   out_data={sign_bit[shift_amt_reg-1:0],in_data[31:shift_amt_reg]};
                  if(shift_amt_reg!=0)
                    carry_out=in_data[shift_amt_reg-1];
                  else
                    carry_out=carry_out;
               end
               
        3'b110 :begin
                if(shift_amt_imm!=0)
                  begin
                    temp=shift_amt_imm;
                    out_data=in_data;
                    while(temp!=0)
                    begin
                      out_data={out_data[0],out_data[31:1]};
                      temp=temp-1;
                    end
               //     out_data={in_data[shift_amt_imm-1:0],in_data[31:shift_amt_imm]};
                    carry_out=in_data[shift_amt_imm-1];
                  end
                else
                 begin
                    carry_out=in_data[0];
                    out_data={carry_in,in_data[31:1]};
                 end
                end
                
        3'b111 :begin
                temp1=shift_amt_reg;
                out_data=in_data;
                while(temp1!=0)
                  begin
                    out_data={out_data[0],out_data[31:1]};
                    temp1=temp1-1;
                  end     //     out_data={in_data[shift_amt_reg-1:0],in_data[31:shift_amt_reg]};
                if(|shift_amt_reg)
                    carry_out=in_data[shift_amt_reg-1];            
                else
                    carry_out=carry_in;
                end
      endcase
    end   // ends if ~imm_or_reg
      else
      out_data=in_data_imm<<2*rotation_code;
    end   //end if enable
    else
      out_data=out_data;
    
  end  //end always block
endmodule
  
